module in_port_test(in_port_num);
	output[31:0] in_port_num;
	assign in_port_num=32'b00110000100100010000001010000011;
 
 
endmodule 